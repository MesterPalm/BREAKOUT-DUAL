
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

-- pMem interface
entity pMem is
  port(
    pAddr : in unsigned(31 downto 0);
    pDataOut : out unsigned(31 downto 0);
    pDataIn : in unsigned(31 downto 0);
    readWrite: in std_logic;
    clk : in std_logic);
end pMem;

architecture Behavioral of pMem is
  
-- program Memory
type p_mem_t is array (0 to 542) of unsigned(31 downto 0);
constant p_mem_c : p_mem_t :=(
--b"0010110111_0010111110_10000_0001_001",
--b"1000100000_0100010110_00000_0001_101",
b"00000_00_0000_0000_00000000000000000",
b"00010_01_0111_0000_00000000000000000",
b"00101_10_1110_0101_11110100000011010",
b"00010_01_1000_0000_00000000000000000",
b"10001_00_0000_1000_10110000000011110",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000010111",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000101000010",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000100000",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000100110",
b"00010_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000111010001",
b"00010_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000001",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000111010001",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000101010",
b"00000_00_0000_0000_00000000000000000",
b"10100_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000010111",
b"10011_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000111",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000101011001",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000010111",
b"10010_01_0111_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"10010_01_1000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000001011",
b"00010_01_0110_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000001101",
b"00101_00_0000_0111_00000000000000000",
b"01111_01_0000_0000_00000000000000000",
b"00000_00_0001_1111_11111000000000000",
b"01011_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"00010_01_0010_0000_00000000000000000",
b"00000_00_0000_0000_00000000000001000",
b"00111_00_0010_0000_00000000000000000",
b"01100_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000010010100",
b"00101_00_0001_0111_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"00101_00_0011_0001_00000000000000000",
b"00101_00_0100_1001_00000000000000000",
b"00111_00_0011_0100_00000000000000000",
b"01100_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000010000110",
b"01101_01_0100_0000_00000000000000000",
b"00000_00_0000_0000_00000000000101110",
b"00111_00_0011_0100_00000000000000000",
b"01100_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000010001010",
b"01101_01_0100_0000_00000000000000000",
b"00000_00_0000_0000_00000000000101110",
b"00111_00_0011_0100_00000000000000000",
b"01100_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000010010000",
b"00010_01_0111_0000_00000000000000000",
b"00101_10_1110_0101_11110100000011010",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000010010100",
b"01111_01_0111_0000_00000000000000000",
b"11111_11_1111_1111_11111111111111000",
b"10000_01_0111_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000101",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000010010100",
b"01111_01_0111_0000_00000000000000000",
b"11111_11_1111_1111_11111111111111000",
b"10000_01_0111_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000111",
b"00010_01_0010_0000_00000000000000000",
b"00000_00_0000_0000_00000000111000000",
b"00111_00_0000_0010_00000000000000000",
b"01100_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000010110101",
b"00101_00_0100_1010_00000000000000000",
b"00111_00_0011_0100_00000000000000000",
b"01100_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000010100111",
b"01101_01_0100_0000_00000000000000000",
b"00000_00_0000_0000_00000000000101110",
b"00111_00_0011_0100_00000000000000000",
b"01100_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000010101011",
b"01101_01_0100_0000_00000000000000000",
b"00000_00_0000_0000_00000000000101110",
b"00111_00_0011_0100_00000000000000000",
b"01100_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000010110001",
b"00010_01_0111_0000_00000000000000000",
b"00101_10_1110_0101_11110100000011010",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000010110101",
b"01111_01_0111_0000_00000000000000000",
b"11111_11_1111_1111_11111111111111000",
b"10000_01_0111_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000011",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000010110101",
b"01111_01_0111_0000_00000000000000000",
b"11111_11_1111_1111_11111111111111000",
b"10000_01_0111_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000001",
b"00101_00_0000_1000_00000000000000000",
b"01111_01_0000_0000_00000000000000000",
b"00000_00_0001_1111_11111000000000000",
b"01011_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"00010_01_0010_0000_00000000000000000",
b"00000_00_0000_0000_00000000000001000",
b"00111_00_0010_0000_00000000000000000",
b"01100_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000100011111",
b"00101_00_0001_1000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01011_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"00101_00_0011_0001_00000000000000000",
b"00101_00_0100_1010_00000000000000000",
b"00111_00_0011_0100_00000000000000000",
b"01100_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000100010001",
b"01101_01_0100_0000_00000000000000000",
b"00000_00_0000_0000_00000000000101110",
b"00111_00_0011_0100_00000000000000000",
b"01100_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000100010101",
b"01101_01_0100_0000_00000000000000000",
b"00000_00_0000_0000_00000000000101110",
b"00111_00_0011_0100_00000000000000000",
b"01100_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000100011011",
b"00010_01_1000_0000_00000000000000000",
b"10001_00_0000_1000_10110000000011110",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000100011111",
b"01111_01_1000_0000_00000000000000000",
b"11111_11_1111_1111_11111111111111000",
b"10000_01_1000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000101",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000100011111",
b"01111_01_1000_0000_00000000000000000",
b"11111_11_1111_1111_11111111111111000",
b"10000_01_1000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000111",
b"00010_01_0010_0000_00000000000000000",
b"00000_00_0000_0000_00000000111010000",
b"00111_00_0000_0010_00000000000000000",
b"01100_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000101000000",
b"00101_00_0100_1010_00000000000000000",
b"00111_00_0011_0100_00000000000000000",
b"01100_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000100110010",
b"01101_01_0100_0000_00000000000000000",
b"00000_00_0000_0000_00000000000101110",
b"00111_00_0011_0100_00000000000000000",
b"01100_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000100110110",
b"01101_01_0100_0000_00000000000000000",
b"00000_00_0000_0000_00000000000101110",
b"00111_00_0011_0100_00000000000000000",
b"01100_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000100111100",
b"00010_01_1000_0000_00000000000000000",
b"10001_00_0000_1000_10110000000011110",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000101000000",
b"01111_01_1000_0000_00000000000000000",
b"11111_11_1111_1111_11111111111111000",
b"10000_01_1000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000011",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000101000000",
b"01111_01_1000_0000_00000000000000000",
b"11111_11_1111_1111_11111111111111000",
b"10000_01_1000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000001",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000010111",
b"00010_01_1111_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000011",
b"00010_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"00010_01_0010_0000_00000000000000000",
b"00000_00_0000_0000_00000000000001111",
b"00010_01_0011_0000_00000000000000000",
b"00000_00_0000_0000_00000000000010010",
b"00010_01_0100_0000_00000000000000000",
b"00000_00_0000_0000_00000000000010011",
b"01000_11_0011_0000_00000001111101000",
b"01101_01_1111_0000_00000000000000000",
b"00000_00_0000_0000_00000000000010000",
b"01000_11_0100_0000_00000001111101000",
b"01101_01_1111_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000100",
b"01101_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000001",
b"00111_00_0001_0010_00000000000000000",
b"00110_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000001001",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000101001100",
b"00010_01_0100_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000011",
b"00111_00_0110_0100_00000000000000000",
b"00110_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000101111000",
b"00101_00_0101_0110_00000000000000000",
b"01111_01_0101_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000001",
b"00010_01_0100_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000001",
b"00111_00_0101_0100_00000000000000000",
b"00110_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000101101011",
b"00010_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000111",
b"00111_00_0000_1011_00000000000000000",
b"01100_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000101111010",
b"00101_00_0101_0110_00000000000000000",
b"01111_01_0101_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000010",
b"00010_01_0100_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000010",
b"00111_00_0101_0100_00000000000000000",
b"00110_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000101111000",
b"00010_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000111",
b"00111_00_0000_1100_00000000000000000",
b"01100_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000110000110",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000011110",
b"00101_00_0001_1011_00000000000000000",
b"01111_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000111",
b"10001_00_0111_0001_00000000000000000",
b"10000_01_0110_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000001",
b"00010_01_0100_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000110010010",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000101101011",
b"00101_00_0010_1100_00000000000000000",
b"01111_01_0010_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000111",
b"10001_00_1000_0010_00000000000000000",
b"10000_01_0110_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000010",
b"00010_01_0100_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000001",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000110010010",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000101111000",
b"00010_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"00111_00_0000_0100_00000000000000000",
b"01001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000110101011",
b"00101_00_1111_1101_00000000000000000",
b"00010_11_0001_0000_00000001111101000",
b"00101_00_0101_0111_00000000000000000",
b"01111_01_0101_0000_00000000000000000",
b"00000_00_0000_0000_00000100000000000",
b"00111_00_0000_0101_00000000000000000",
b"00110_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000110100101",
b"00010_10_0010_0000_00000000111001111",
b"01101_01_0010_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000001",
b"01000_10_0010_0000_00000000111001111",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000110111101",
b"00010_10_0010_0000_00000000111010000",
b"01101_01_0010_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000001",
b"01000_10_0010_0000_00000000111010000",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000110111101",
b"00101_00_1111_1110_00000000000000000",
b"00010_11_0001_0000_00000001111101000",
b"00101_00_0101_1000_00000000000000000",
b"01111_01_0101_0000_00000000000000000",
b"00000_00_0000_0000_00000100000000000",
b"00111_00_0000_0101_00000000000000000",
b"00110_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000110111001",
b"00010_10_0010_0000_00000000111001111",
b"01101_01_0010_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000001",
b"01000_10_0010_0000_00000000111001111",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000110111101",
b"00010_10_0010_0000_00000000111010000",
b"01101_01_0010_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000001",
b"01000_10_0010_0000_00000000111010000",
b"00010_01_0010_0000_00000000000000000",
b"00000_00_0000_0000_00000000000010010",
b"00111_00_0001_0010_00000000000000000",
b"00110_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000111001010",
b"00010_01_0010_0000_00000000000000000",
b"00000_00_0000_0000_00000000000010011",
b"00111_00_0001_0010_00000000000000000",
b"00110_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000111001010",
b"00010_01_0101_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01000_11_0101_0000_00000001111101000",
b"00111_00_0000_0100_00000000000000000",
b"00110_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000110000100",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000110010000",
b"00000_00_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"00010_01_0010_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"00111_00_0001_0010_00000000000000000",
b"00110_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000111011011",
b"00010_10_0011_0000_00000000111010000",
b"00010_01_1111_0000_00000000000000000",
b"00000_00_0000_0000_00000000100011000",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000111011110",
b"00010_10_0011_0000_00000000111001111",
b"00010_01_1111_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01110_01_0011_0000_00000000000000000",
b"00000_00_0000_0000_00000000001100100",
b"01100_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000111100110",
b"01101_01_0010_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000001",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000111011110",
b"01101_01_0011_0000_00000000000000000",
b"00000_00_0000_0000_00000000001100100",
b"00010_01_0100_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"00111_00_0010_0100_00000000000000000",
b"01001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000111101111",
b"00010_01_0010_0000_00000000000000000",
b"00000_00_0000_0000_00000000000001010",
b"01000_11_0010_0000_00000001111101000",
b"00010_01_0010_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01110_01_0011_0000_00000000000000000",
b"00000_00_0000_0000_00000000000001010",
b"01100_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000111111010",
b"01101_01_0010_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000001",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000111110010",
b"01101_01_0011_0000_00000000000000000",
b"00000_00_0000_0000_00000000000001010",
b"00111_00_0010_0100_00000000000000000",
b"01001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000001000000001",
b"00010_01_0010_0000_00000000000000000",
b"00000_00_0000_0000_00000000000001010",
b"01101_01_1111_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000001",
b"01000_11_0010_0000_00000001111101000",
b"00010_01_0010_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"01110_01_0011_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000001",
b"01100_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000001000001110",
b"01101_01_0010_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000001",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000001000000110",
b"01101_01_0011_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000001",
b"00111_00_0010_0100_00000000000000000",
b"01001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000001000010101",
b"00010_01_0010_0000_00000000000000000",
b"00000_00_0000_0000_00000000000001010",
b"01101_01_1111_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000001",
b"01000_11_0010_0000_00000001111101000",
b"00010_01_0010_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"00111_00_0001_0010_00000000000000000",
b"00110_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000010001",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000010101"
);

   signal p_mem : p_mem_t := p_mem_c;

begin  -- pMem
  -- purpose: data in or data out 
  pDataOut <= p_mem(to_integer(pAddr)) when (readWrite = '1') else
                    (others => '0');
  
  process (clk)
  begin  -- process
    if(rising_edge(clk)) then
      if (readWrite = '0') then
        p_mem(to_integer(pAddr)) <= pDataIn;
      end if;
    end if;       
  end process;
 
end Behavioral;
