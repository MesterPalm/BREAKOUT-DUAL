
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

-- pMem interface
entity pMem is
  port(
    pAddr : in unsigned(31 downto 0);
    pDataOut : out unsigned(31 downto 0);
    pDataIn : in unsigned(31 downto 0);
    readWrite: in std_logic;
    clk : in std_logic);
end pMem;

architecture Behavioral of pMem is

-- program Memory
type p_mem_t is array (0 to 44) of unsigned(31 downto 0);
constant p_mem_c : p_mem_t :=(
b"00000_00_0000_0000_00000000000000000",
b"00010_01_0111_0000_00000000000000000",
b"01000_00_1000_1110_00000000000001001",
b"00010_01_1000_0000_00000000000000000",
b"01100_00_0000_1110_00000000000001001",--------------------------
b"00010_01_1111_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"00010_01_0110_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"00010_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000001000",
b"00010_01_0110_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000001",
b"00010_01_0110_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"10010_01_0111_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"10010_01_1000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000000",
b"00111_00_0000_1011_00000000000000000",
b"01100_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000011011",
b"00111_00_0000_1100_00000000000000000",
b"01100_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000100010",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000100111",
b"00101_00_0001_1011_00000000000000000",
b"01111_01_0001_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000111",
b"01000_11_0001_0000_00000001111101000",
b"10001_00_0111_0001_00000000000000000",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000010110",
b"00101_00_0010_1100_00000000000000000",
b"01111_01_0010_0000_00000000000000000",
b"00000_00_0000_0000_00000000000000111",
b"01000_11_0010_0000_00000001111101001",
b"10001_00_1000_0010_00000000000000000",
b"10011_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000001111",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000010011",
b"00001_01_0000_0000_00000000000000000",
b"00000_00_0000_0000_00000000000100111"


);

   signal p_mem : p_mem_t := p_mem_c;

begin  -- pMem
  -- purpose: data in or data out 
  pDataOut <= p_mem(to_integer(pAddr)) when (readWrite = '1') else
                    (others => '0');
  
  process (clk)
  begin  -- process
    if(rising_edge(clk)) then
      if (readWrite = '0') then
        p_mem(to_integer(pAddr)) <= pDataIn;
      end if;
    end if;       
  end process;
 
end Behavioral;
