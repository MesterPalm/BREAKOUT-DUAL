
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

-- pMem interface
entity pMem is
  port(
    pAddr : in unsigned(31 downto 0);
    pDataOut : out unsigned(31 downto 0);
    pDataIn : in unsigned(31 downto 0);
    readWrite: in std_logic;
    clk : in std_logic);
end pMem;

architecture Behavioral of pMem is

-- program Memory
type p_mem_t is array (0 to 451) of unsigned(31 downto 0);
constant p_mem_c : p_mem_t :=(
  b"00000_00_0000_0000_00000000000000000",
  b"00010_01_0111_0000_00000000000000000",
  b"00000_00_0000_0011_00000000000000110",
  b"00010_01_1000_0000_00000000000000000",
  b"00000_00_0000_0111_00000000000000010",
  b"00001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000010001",
  b"00001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000010101",
  b"00010_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"00001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000101110100",
  b"00010_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000001",
  b"00001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000101110100",
  b"10011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000111",
  b"00001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000010001",
  b"10010_01_0111_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"10010_01_1000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"00001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000001001",
  b"00010_01_0110_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"00001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000001001",
  b"00101_00_0000_0111_00000000000000000",
  b"01111_01_0000_0000_00000000000000000",
  b"00000_00_0000_1111_11111000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"00010_01_0010_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000001000",
  b"00111_00_0000_0010_00000000000000000",
  b"01100_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000010000111",
  b"00101_00_0001_0111_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"00101_00_0011_0001_00000000000000000",
  b"00101_00_0100_1001_00000000000000000",
  b"00111_00_0011_0100_00000000000000000",
  b"01100_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000010000111",
  b"01101_01_0100_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000101110",
  b"00111_00_0011_0100_00000000000000000",
  b"01100_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000100010000",
  b"01101_01_0100_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000101110",
  b"00111_00_0011_0100_00000000000000000",
  b"01100_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000100010110",
  b"00001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000010000111",
  b"01111_01_0111_0000_00000000000000000",
  b"00000_00_0000_1111_11111111111111000",
  b"10000_01_0111_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000101",
  b"00001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000010000111",
  b"01111_01_0111_0000_00000000000000000",
  b"00000_00_0000_1111_11111111111111000",
  b"10000_01_0111_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000111",
  b"00010_01_0010_0000_00000000000000000",
  b"00000_00_0000_0000_00000000111011000",
  b"00111_00_0000_0010_00000000000000000",
  b"01100_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000010100110",
  b"00101_00_0100_1010_00000000000000000",
  b"00111_00_0011_0100_00000000000000000",
  b"01100_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000010100110",
  b"01101_01_0100_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000101110",
  b"00111_00_0011_0100_00000000000000000",
  b"01100_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000100101111",
  b"01101_01_0100_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000101110",
  b"00111_00_0011_0100_00000000000000000",
  b"01100_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000100110101",
  b"00001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000010100110",
  b"01111_01_0111_0000_00000000000000000",
  b"00000_00_0000_1111_11111111111111000",
  b"10000_01_0111_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000011",
  b"00001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000010100110",
  b"01111_01_0111_0000_00000000000000000",
  b"00000_00_0000_1111_11111111111111000",
  b"10000_01_0111_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000001",
  b"00101_00_0000_1000_00000000000000000",
  b"01111_01_0000_0000_00000000000000000",
  b"00000_00_0000_1111_11111000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"00010_01_0010_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000001000",
  b"00111_00_0000_0010_00000000000000000",
  b"01100_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000100011010",
  b"00101_00_0001_1000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01011_01_0001_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"00101_00_0011_0000_00000000000000000",
  b"00101_00_0100_1001_00000000000000000",
  b"00111_00_0011_0100_00000000000000000",
  b"01100_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000100011010",
  b"01101_01_0100_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000101110",
  b"00111_00_0011_0100_00000000000000000",
  b"01100_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000001111101",
  b"01101_01_0100_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000101110",
  b"00111_00_0011_0100_00000000000000000",
  b"01100_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000010000011",
  b"00001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000100011010",
  b"01111_01_1000_0000_00000000000000000",
  b"00000_00_0000_1111_11111111111111000",
  b"10000_01_1000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000101",
  b"00001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000100011010",
  b"01111_01_1000_0000_00000000000000000",
  b"00000_00_0000_1111_11111111111111000",
  b"10000_01_1000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000111",
  b"00010_01_0010_0000_00000000000000000",
  b"00000_00_0000_0000_00000000111011000",
  b"00111_00_0000_0010_00000000000000000",
  b"01100_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000100111001",
  b"00101_00_0100_1010_00000000000000000",
  b"00111_00_0011_0100_00000000000000000",
  b"01100_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000100111001",
  b"01101_01_0100_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000101110",
  b"00111_00_0011_0100_00000000000000000",
  b"01100_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000010011100",
  b"01101_01_0100_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000101110",
  b"00111_00_0011_0100_00000000000000000",
  b"01100_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000010100010",
  b"00001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000100111001",
  b"01111_01_1000_0000_00000000000000000",
  b"00000_00_0000_1111_11111111111111000",
  b"10000_01_1000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000011",
  b"00001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000100111001",
  b"01111_01_1000_0000_00000000000000000",
  b"00000_00_0000_1111_11111111111111000",
  b"10000_01_1000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000001",
  b"00001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000010011",
  b"00010_01_0101_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000011",
  b"00111_00_0110_0101_00000000000000000",
  b"00110_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000101100001",
  b"00010_01_0101_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000001",
  b"00111_00_0110_0101_00000000000000000",
  b"00110_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000101010011",
  b"00010_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000001000",
  b"00111_00_1011_0000_00000000000000000",
  b"01100_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000101010011",
  b"00101_00_0011_1011_00000000000000000",
  b"01111_01_0011_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000111",
  b"10001_00_0111_0011_00000000000000000",
  b"01101_01_0110_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000001",
  b"00101_00_0000_1101_00000000000000000",
  b"00001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000101100011",
  b"00010_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000001000",
  b"00111_00_1100_0000_00000000000000000",
  b"01100_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000101100001",
  b"00101_00_0100_1100_00000000000000000",
  b"01111_01_0100_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000111",
  b"10001_00_1000_0100_00000000000000000",
  b"01101_01_0110_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000010",
  b"00101_00_0000_1101_00000000000000000",
  b"00001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000101100011",
  b"00001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000010011",
  b"00101_00_1111_0000_00000000000000000",
  b"00010_11_0001_0000_00000001111101000",
  b"00010_01_0010_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000010010",
  b"00111_00_0001_0010_00000000000000000",
  b"00110_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000101110010",
  b"00010_01_0010_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000010011",
  b"00111_00_0001_0010_00000000000000000",
  b"00110_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000101110010",
  b"00010_01_0011_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01000_11_0011_0000_00000001111101000",
  b"00001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000010001",
  b"00000_00_0000_0000_00000000001100100",
  b"00000_00_0000_0000_00000000001100100",
  b"00010_01_0010_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"00111_00_0001_0010_00000000000000000",
  b"00110_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000101111110",
  b"00010_10_0011_0000_00000000101110101",
  b"00010_01_1111_0000_00000000000000000",
  b"00000_00_0000_0000_00000000100011000",
  b"00001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000110000001",
  b"00010_10_0011_0000_00000000101110100",
  b"00010_01_1111_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01110_01_0011_0000_00000000000000000",
  b"00000_00_0000_0000_00000000001100100",
  b"01100_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000110001001",
  b"01101_01_0010_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000001",
  b"00001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000110000011",
  b"01101_01_0011_0000_00000000000000000",
  b"00000_00_0000_0000_00000000001100100",
  b"00010_01_0100_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"00111_00_0010_0100_00000000000000000",
  b"01001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000110010010",
  b"00010_01_0010_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000001010",
  b"01000_11_0010_0000_00000001111101000",
  b"00010_01_0010_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01110_01_0011_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000001010",
  b"01100_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000110011101",
  b"01101_01_0010_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000001",
  b"00001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000110010111",
  b"01101_01_0011_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000001010",
  b"00111_00_0010_0100_00000000000000000",
  b"01001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000110100100",
  b"00010_01_0010_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000001010",
  b"01101_01_1111_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000001",
  b"01000_11_0010_0000_00000001111101000",
  b"00010_01_0010_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"01110_01_0011_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000001",
  b"01100_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000110110001",
  b"01101_01_0010_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000001",
  b"00001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000110101011",
  b"01101_01_0011_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000001",
  b"00111_00_0010_0100_00000000000000000",
  b"01001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000110111000",
  b"00010_01_0010_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000001010",
  b"01101_01_1111_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000001",
  b"01000_11_0010_0000_00000001111101000",
  b"00010_01_0010_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000000000",
  b"00111_00_0001_0010_00000000000000000",
  b"00110_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000001101",
  b"00001_01_0000_0000_00000000000000000",
  b"00000_00_0000_0000_00000000000010001");

   signal p_mem : p_mem_t := p_mem_c;

begin  -- pMem
  -- purpose: data in or data out 
  pDataOut <= p_mem(to_integer(pAddr)) when (readWrite = '1') else
                    (others => '0');
  
  process (clk)
  begin  -- process
    if(rising_edge(clk)) then
      if (readWrite = '1') then
        p_mem(to_integer(pAddr)) <= pDataIn;
      end if;
    end if;       
  end process;
 
end Behavioral;
