
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

-- pMem interface
entity pMem is
  port(
    pAddr : in unsigned(31 downto 0);
    pDataOut : out unsigned(31 downto 0);
    pDataIn : in unsigned(31 downto 0);
    readWrite: in std_logic);
end pMem;

architecture Behavioral of pMem is

-- program Memory
type p_mem_t is array (0 to 11) of unsigned(31 downto 0);
constant p_mem_c : p_mem_t :=
--(X"12200000",
-- X"000000C4",
-- X"12400000",
-- X"00000001",
-- X"18420000");
   --(b"00010_01_0001_0000_00000000000000000",  --0 LOAD GR 0001 0111          
   -- b"00000_00_0000_0000_00000000000001110",  --1  
   -- b"00010_01_0010_0000_00000000000000000",  --10  LOAD GR 0010 0001
   -- b"00000_00_0000000000000000000000001",  --11        
   -- b"00010_01_0011_0000_00000000000000000",  --100 LOAD GR 0011 0001 
   -- b"00000_00_0000_0000_00000000000000001",  --101
   -- b"00011_00_0011_0010_00000000000000000",  --110 ADD GR 0011 GR 0010        
   -- b"00111_00_0011_0001_00000000000000000",  --111 CMP GR 0011 GR 0111
   -- b"00110_01_0000_0000_00000000000000000", --1000 BEQ  1011
   -- b"00000_00_0000000000000000000001111",  --1001    
   -- b"00001_01_0000000000000000000000000",  --1010   BRA 
   -- b"00000_00_0000000000000000000000110",  --1011
   -- b"00000_00_0000000000000000000000000",  --1100
   -- b"00000_00_0000000000000000000000000",  --1101
   -- b"00000_00_0000000000000000000000000",  --1110   
   -- b"00000_00_0000000000000000000000000"); --1111
  --(b"00000_00_0000000000000000000000000",
  --  b"00010_01_0001_000000000000000000000",
  -- b"00001_01_0000000000000000000000000",
  -- b"01000_10_0001_000000000000000001110",
  -- b"00000_00_0000000000000000000000000",
  -- b"00000_00_0000000000000000000000000",
  -- b"00000_00_0000000000000000000000000",
  -- b"00000_00_0000000000000000000000000",
  -- b"00000_00_0000000000000000000000000",
  -- b"00000_00_0000000000000000000000000",
  -- b"00000_00_0000000000000000000000000",
  -- b"00000_00_0000000000000000000000000",
  -- b"00000_00_0000000000000000000000000",
  -- b"00000_00_0000000000000000000000000",
  -- b"00000_00_0000000000000000000000000",
  -- b"00000_00_0000000000000000000000001");
  (b"00010_01_0010_0000_00000000000000000",
   b"00000_00_0000_0000_00000000000000111",
   b"00010_01_0011_0000_00000000000000000",
   b"10000_00_0000_0000_00000000000011111",
   b"01011_00_0011_0000_00000000000000000",
   b"00001_01_0000_0000_00000000000000000",
   b"00000_00_0000_0000_00000000000000100",
   b"00000_00_0000_0000_00000000000000000",
   b"00000_00_0000_0000_00000000000000000",
   b"00000_00_0000_0000_00000000000000000",
   b"00000_00_0000_0000_00000000000000000",
   b"00000_00_0000_0000_00000000000000000"
   );

   signal p_mem : p_mem_t := p_mem_c;

begin  -- pMem
  -- purpose: data in or data out 
  process (readWrite, pAddr)
  begin  -- process
    if (readWrite = '1') then
       pDataOut <= p_mem(to_integer(pAddr));
    elsif (readWrite = '0') then
      p_mem(to_integer(pAddr)) <= pDataIn;
    end if;
  end process;
 
end Behavioral;
