library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

-- pMem interface
entity pMem is
  port(
    pAddr : in unsigned(31 downto 0);
    pData : out unsigned(31 downto 0));
end pMem;

architecture Behavioral of pMem is

-- program Memory
type p_mem_t is array (0 to 15) of unsigned(31 downto 0);
constant p_mem_c : p_mem_t :=
  (b"00010_01_0001_0000_00000000000000000",  --0 LOAD GR 0001 0111          
   b"00000_00_0000_0000_00000000000000010",  --1  
   b"00010_01_0010_0000_00000000000000000",  --10  LOAD GR 0010 0001
   b"00000_00_0000000000000000000000001",  --11        
   b"00010_01_0011_0000_00000000000000000",  --100 LOAD GR 0011 0001 
   b"00000_00_0000_0000_00000000000000001",  --101
   b"00011_00_0011_0010_00000000000000000",  --110 ADD GR 0011 GR 0010        
   b"00111_00_0011_0001_00000000000000000",  --111 CMP GR 0011 GR 0111
   b"00110_01_0000_0000_00000000000000000", --1000 BEQ  1011
   b"00000_00_0000000000000000000001111",  --1001    
   b"00001_01_0000000000000000000000000",  --1010   BRA 
   b"00000_00_0000000000000000000000000",  --1011
   b"00000_00_0000000000000000000000000",  --1100
   b"00000_00_0000000000000000000000000",  --1101
   b"00000_00_0000000000000000000000000",  --1110   
   b"00000_00_0000000000000000000000000"); --1111

  signal p_mem : p_mem_t := p_mem_c;


begin  -- pMem
  pData <= p_mem(to_integer(pAddr));

end Behavioral;
